module test();
	wire[15:0]x;
	wire[9:0]y = 10'b0001110001;
	assign x = y;
endmodule
